//`timescale 1ns / 1ps
module me_sad_calculation (clk, search, current, SAD01, SAD02, SAD03, SAD04, SAD05, SAD06, SAD07, SAD08, SAD09, SAD10, SAD11, SAD12, SAD13, SAD14, SAD15, SAD16);
	
	input clk;
	
	input [((8*16*17)-1):0] search;
	input [((8*16*16)-1):0] current;
	output reg [11:0] SAD01, SAD02, SAD03, SAD04, SAD05, SAD06, SAD07, SAD08, SAD09, SAD10, SAD11, SAD12, SAD13, SAD14, SAD15, SAD16;
		
	wire [7:0] difference_matrix [15:0][15:0];
	
	reg [9:0] add01, add02, add03, add04, add05, add06, add07, add08, add09, add10, add11, add12, add13, add14, add15, add16, add17, add18, add19, add20, add21, add22, add23, add24, add25, add26, add27, add28, add29, add30, add31, add32;
	reg [9:0] add33, add34, add35, add36, add37, add38, add39, add40, add41, add42, add43, add44, add45, add46, add47, add48, add49, add50, add51, add52, add53, add54, add55, add56, add57, add58, add59, add60, add61, add62, add63, add64;

me_PE PE_ij256 (.clk(clk),.A(search[((8*((17*0)+0 +2))-1):(8*((17*0)+0 +1))]),.B(current[((8*((16*0)+0 +1))-1):(8*((16*0)+0 ))]),.AD(difference_matrix[0][0 ]));
me_PE PE_ij241 (.clk(clk),.A(search[((8*((17*0)+1 +2))-1):(8*((17*0)+1 +1))]),.B(current[((8*((16*0)+1 +1))-1):(8*((16*0)+1 ))]),.AD(difference_matrix[0][1 ]));
me_PE PE_ij242 (.clk(clk),.A(search[((8*((17*0)+2 +2))-1):(8*((17*0)+2 +1))]),.B(current[((8*((16*0)+2 +1))-1):(8*((16*0)+2 ))]),.AD(difference_matrix[0][2 ]));
me_PE PE_ij243 (.clk(clk),.A(search[((8*((17*0)+3 +2))-1):(8*((17*0)+3 +1))]),.B(current[((8*((16*0)+3 +1))-1):(8*((16*0)+3 ))]),.AD(difference_matrix[0][3 ]));
me_PE PE_ij244 (.clk(clk),.A(search[((8*((17*0)+4 +2))-1):(8*((17*0)+4 +1))]),.B(current[((8*((16*0)+4 +1))-1):(8*((16*0)+4 ))]),.AD(difference_matrix[0][4 ]));
me_PE PE_ij245 (.clk(clk),.A(search[((8*((17*0)+5 +2))-1):(8*((17*0)+5 +1))]),.B(current[((8*((16*0)+5 +1))-1):(8*((16*0)+5 ))]),.AD(difference_matrix[0][5 ]));
me_PE PE_ij246 (.clk(clk),.A(search[((8*((17*0)+6 +2))-1):(8*((17*0)+6 +1))]),.B(current[((8*((16*0)+6 +1))-1):(8*((16*0)+6 ))]),.AD(difference_matrix[0][6 ]));
me_PE PE_ij247 (.clk(clk),.A(search[((8*((17*0)+7 +2))-1):(8*((17*0)+7 +1))]),.B(current[((8*((16*0)+7 +1))-1):(8*((16*0)+7 ))]),.AD(difference_matrix[0][7 ]));
me_PE PE_ij248 (.clk(clk),.A(search[((8*((17*0)+8 +2))-1):(8*((17*0)+8 +1))]),.B(current[((8*((16*0)+8 +1))-1):(8*((16*0)+8 ))]),.AD(difference_matrix[0][8 ]));
me_PE PE_ij249 (.clk(clk),.A(search[((8*((17*0)+9 +2))-1):(8*((17*0)+9 +1))]),.B(current[((8*((16*0)+9 +1))-1):(8*((16*0)+9 ))]),.AD(difference_matrix[0][9 ]));
me_PE PE_ij250 (.clk(clk),.A(search[((8*((17*0)+10+2))-1):(8*((17*0)+10+1))]),.B(current[((8*((16*0)+10+1))-1):(8*((16*0)+10))]),.AD(difference_matrix[0][10]));
me_PE PE_ij251 (.clk(clk),.A(search[((8*((17*0)+11+2))-1):(8*((17*0)+11+1))]),.B(current[((8*((16*0)+11+1))-1):(8*((16*0)+11))]),.AD(difference_matrix[0][11]));
me_PE PE_ij252 (.clk(clk),.A(search[((8*((17*0)+12+2))-1):(8*((17*0)+12+1))]),.B(current[((8*((16*0)+12+1))-1):(8*((16*0)+12))]),.AD(difference_matrix[0][12]));
me_PE PE_ij253 (.clk(clk),.A(search[((8*((17*0)+13+2))-1):(8*((17*0)+13+1))]),.B(current[((8*((16*0)+13+1))-1):(8*((16*0)+13))]),.AD(difference_matrix[0][13]));
me_PE PE_ij254 (.clk(clk),.A(search[((8*((17*0)+14+2))-1):(8*((17*0)+14+1))]),.B(current[((8*((16*0)+14+1))-1):(8*((16*0)+14))]),.AD(difference_matrix[0][14]));
me_PE PE_ij255 (.clk(clk),.A(search[((8*((17*0)+15+2))-1):(8*((17*0)+15+1))]),.B(current[((8*((16*0)+15+1))-1):(8*((16*0)+15))]),.AD(difference_matrix[0][15]));
	
	
me_PE PE_ij16 (.clk(clk),.A(search[((8*((17*1)+0 +2))-1):(8*((17*1)+0 +1))]),.B(current[((8*((16*1)+0 +1))-1):(8*((16*1)+0 ))]),.AD(difference_matrix[1][0 ]));
me_PE PE_ij1  (.clk(clk),.A(search[((8*((17*1)+1 +2))-1):(8*((17*1)+1 +1))]),.B(current[((8*((16*1)+1 +1))-1):(8*((16*1)+1 ))]),.AD(difference_matrix[1][1 ]));
me_PE PE_ij2  (.clk(clk),.A(search[((8*((17*1)+2 +2))-1):(8*((17*1)+2 +1))]),.B(current[((8*((16*1)+2 +1))-1):(8*((16*1)+2 ))]),.AD(difference_matrix[1][2 ]));
me_PE PE_ij3  (.clk(clk),.A(search[((8*((17*1)+3 +2))-1):(8*((17*1)+3 +1))]),.B(current[((8*((16*1)+3 +1))-1):(8*((16*1)+3 ))]),.AD(difference_matrix[1][3 ]));
me_PE PE_ij4  (.clk(clk),.A(search[((8*((17*1)+4 +2))-1):(8*((17*1)+4 +1))]),.B(current[((8*((16*1)+4 +1))-1):(8*((16*1)+4 ))]),.AD(difference_matrix[1][4 ]));
me_PE PE_ij5  (.clk(clk),.A(search[((8*((17*1)+5 +2))-1):(8*((17*1)+5 +1))]),.B(current[((8*((16*1)+5 +1))-1):(8*((16*1)+5 ))]),.AD(difference_matrix[1][5 ]));
me_PE PE_ij6  (.clk(clk),.A(search[((8*((17*1)+6 +2))-1):(8*((17*1)+6 +1))]),.B(current[((8*((16*1)+6 +1))-1):(8*((16*1)+6 ))]),.AD(difference_matrix[1][6 ]));
me_PE PE_ij7  (.clk(clk),.A(search[((8*((17*1)+7 +2))-1):(8*((17*1)+7 +1))]),.B(current[((8*((16*1)+7 +1))-1):(8*((16*1)+7 ))]),.AD(difference_matrix[1][7 ]));
me_PE PE_ij8  (.clk(clk),.A(search[((8*((17*1)+8 +2))-1):(8*((17*1)+8 +1))]),.B(current[((8*((16*1)+8 +1))-1):(8*((16*1)+8 ))]),.AD(difference_matrix[1][8 ]));
me_PE PE_ij9  (.clk(clk),.A(search[((8*((17*1)+9 +2))-1):(8*((17*1)+9 +1))]),.B(current[((8*((16*1)+9 +1))-1):(8*((16*1)+9 ))]),.AD(difference_matrix[1][9 ]));
me_PE PE_ij10 (.clk(clk),.A(search[((8*((17*1)+10+2))-1):(8*((17*1)+10+1))]),.B(current[((8*((16*1)+10+1))-1):(8*((16*1)+10))]),.AD(difference_matrix[1][10]));
me_PE PE_ij11 (.clk(clk),.A(search[((8*((17*1)+11+2))-1):(8*((17*1)+11+1))]),.B(current[((8*((16*1)+11+1))-1):(8*((16*1)+11))]),.AD(difference_matrix[1][11]));
me_PE PE_ij12 (.clk(clk),.A(search[((8*((17*1)+12+2))-1):(8*((17*1)+12+1))]),.B(current[((8*((16*1)+12+1))-1):(8*((16*1)+12))]),.AD(difference_matrix[1][12]));
me_PE PE_ij13 (.clk(clk),.A(search[((8*((17*1)+13+2))-1):(8*((17*1)+13+1))]),.B(current[((8*((16*1)+13+1))-1):(8*((16*1)+13))]),.AD(difference_matrix[1][13]));
me_PE PE_ij14 (.clk(clk),.A(search[((8*((17*1)+14+2))-1):(8*((17*1)+14+1))]),.B(current[((8*((16*1)+14+1))-1):(8*((16*1)+14))]),.AD(difference_matrix[1][14]));
me_PE PE_ij15 (.clk(clk),.A(search[((8*((17*1)+15+2))-1):(8*((17*1)+15+1))]),.B(current[((8*((16*1)+15+1))-1):(8*((16*1)+15))]),.AD(difference_matrix[1][15]));


me_PE PE_ij32 (.clk(clk),.A(search[((8*((17*2)+0 +2))-1):(8*((17*2)+0 +1))]),.B(current[((8*((16*2)+0 +1))-1):(8*((16*2)+0 ))]),.AD(difference_matrix[2][0 ]));
me_PE PE_ij17 (.clk(clk),.A(search[((8*((17*2)+1 +2))-1):(8*((17*2)+1 +1))]),.B(current[((8*((16*2)+1 +1))-1):(8*((16*2)+1 ))]),.AD(difference_matrix[2][1 ]));
me_PE PE_ij18 (.clk(clk),.A(search[((8*((17*2)+2 +2))-1):(8*((17*2)+2 +1))]),.B(current[((8*((16*2)+2 +1))-1):(8*((16*2)+2 ))]),.AD(difference_matrix[2][2 ]));
me_PE PE_ij19 (.clk(clk),.A(search[((8*((17*2)+3 +2))-1):(8*((17*2)+3 +1))]),.B(current[((8*((16*2)+3 +1))-1):(8*((16*2)+3 ))]),.AD(difference_matrix[2][3 ]));
me_PE PE_ij20 (.clk(clk),.A(search[((8*((17*2)+4 +2))-1):(8*((17*2)+4 +1))]),.B(current[((8*((16*2)+4 +1))-1):(8*((16*2)+4 ))]),.AD(difference_matrix[2][4 ]));
me_PE PE_ij21 (.clk(clk),.A(search[((8*((17*2)+5 +2))-1):(8*((17*2)+5 +1))]),.B(current[((8*((16*2)+5 +1))-1):(8*((16*2)+5 ))]),.AD(difference_matrix[2][5 ]));
me_PE PE_ij22 (.clk(clk),.A(search[((8*((17*2)+6 +2))-1):(8*((17*2)+6 +1))]),.B(current[((8*((16*2)+6 +1))-1):(8*((16*2)+6 ))]),.AD(difference_matrix[2][6 ]));
me_PE PE_ij23 (.clk(clk),.A(search[((8*((17*2)+7 +2))-1):(8*((17*2)+7 +1))]),.B(current[((8*((16*2)+7 +1))-1):(8*((16*2)+7 ))]),.AD(difference_matrix[2][7 ]));
me_PE PE_ij24 (.clk(clk),.A(search[((8*((17*2)+8 +2))-1):(8*((17*2)+8 +1))]),.B(current[((8*((16*2)+8 +1))-1):(8*((16*2)+8 ))]),.AD(difference_matrix[2][8 ]));
me_PE PE_ij25 (.clk(clk),.A(search[((8*((17*2)+9 +2))-1):(8*((17*2)+9 +1))]),.B(current[((8*((16*2)+9 +1))-1):(8*((16*2)+9 ))]),.AD(difference_matrix[2][9 ]));
me_PE PE_ij26 (.clk(clk),.A(search[((8*((17*2)+10+2))-1):(8*((17*2)+10+1))]),.B(current[((8*((16*2)+10+1))-1):(8*((16*2)+10))]),.AD(difference_matrix[2][10]));
me_PE PE_ij27 (.clk(clk),.A(search[((8*((17*2)+11+2))-1):(8*((17*2)+11+1))]),.B(current[((8*((16*2)+11+1))-1):(8*((16*2)+11))]),.AD(difference_matrix[2][11]));
me_PE PE_ij28 (.clk(clk),.A(search[((8*((17*2)+12+2))-1):(8*((17*2)+12+1))]),.B(current[((8*((16*2)+12+1))-1):(8*((16*2)+12))]),.AD(difference_matrix[2][12]));
me_PE PE_ij29 (.clk(clk),.A(search[((8*((17*2)+13+2))-1):(8*((17*2)+13+1))]),.B(current[((8*((16*2)+13+1))-1):(8*((16*2)+13))]),.AD(difference_matrix[2][13]));
me_PE PE_ij30 (.clk(clk),.A(search[((8*((17*2)+14+2))-1):(8*((17*2)+14+1))]),.B(current[((8*((16*2)+14+1))-1):(8*((16*2)+14))]),.AD(difference_matrix[2][14]));
me_PE PE_ij31 (.clk(clk),.A(search[((8*((17*2)+15+2))-1):(8*((17*2)+15+1))]),.B(current[((8*((16*2)+15+1))-1):(8*((16*2)+15))]),.AD(difference_matrix[2][15]));

me_PE PE_ij48 (.clk(clk),.A(search[((8*((17*3)+0 +2))-1):(8*((17*3)+0 +1))]),.B(current[((8*((16*3)+0 +1))-1):(8*((16*3)+0 ))]),.AD(difference_matrix[3][0 ]));
me_PE PE_ij33 (.clk(clk),.A(search[((8*((17*3)+1 +2))-1):(8*((17*3)+1 +1))]),.B(current[((8*((16*3)+1 +1))-1):(8*((16*3)+1 ))]),.AD(difference_matrix[3][1 ]));
me_PE PE_ij34 (.clk(clk),.A(search[((8*((17*3)+2 +2))-1):(8*((17*3)+2 +1))]),.B(current[((8*((16*3)+2 +1))-1):(8*((16*3)+2 ))]),.AD(difference_matrix[3][2 ]));
me_PE PE_ij35 (.clk(clk),.A(search[((8*((17*3)+3 +2))-1):(8*((17*3)+3 +1))]),.B(current[((8*((16*3)+3 +1))-1):(8*((16*3)+3 ))]),.AD(difference_matrix[3][3 ]));
me_PE PE_ij36 (.clk(clk),.A(search[((8*((17*3)+4 +2))-1):(8*((17*3)+4 +1))]),.B(current[((8*((16*3)+4 +1))-1):(8*((16*3)+4 ))]),.AD(difference_matrix[3][4 ]));
me_PE PE_ij37 (.clk(clk),.A(search[((8*((17*3)+5 +2))-1):(8*((17*3)+5 +1))]),.B(current[((8*((16*3)+5 +1))-1):(8*((16*3)+5 ))]),.AD(difference_matrix[3][5 ]));
me_PE PE_ij38 (.clk(clk),.A(search[((8*((17*3)+6 +2))-1):(8*((17*3)+6 +1))]),.B(current[((8*((16*3)+6 +1))-1):(8*((16*3)+6 ))]),.AD(difference_matrix[3][6 ]));
me_PE PE_ij39 (.clk(clk),.A(search[((8*((17*3)+7 +2))-1):(8*((17*3)+7 +1))]),.B(current[((8*((16*3)+7 +1))-1):(8*((16*3)+7 ))]),.AD(difference_matrix[3][7 ]));
me_PE PE_ij40 (.clk(clk),.A(search[((8*((17*3)+8 +2))-1):(8*((17*3)+8 +1))]),.B(current[((8*((16*3)+8 +1))-1):(8*((16*3)+8 ))]),.AD(difference_matrix[3][8 ]));
me_PE PE_ij41 (.clk(clk),.A(search[((8*((17*3)+9 +2))-1):(8*((17*3)+9 +1))]),.B(current[((8*((16*3)+9 +1))-1):(8*((16*3)+9 ))]),.AD(difference_matrix[3][9 ]));
me_PE PE_ij42 (.clk(clk),.A(search[((8*((17*3)+10+2))-1):(8*((17*3)+10+1))]),.B(current[((8*((16*3)+10+1))-1):(8*((16*3)+10))]),.AD(difference_matrix[3][10]));
me_PE PE_ij43 (.clk(clk),.A(search[((8*((17*3)+11+2))-1):(8*((17*3)+11+1))]),.B(current[((8*((16*3)+11+1))-1):(8*((16*3)+11))]),.AD(difference_matrix[3][11]));
me_PE PE_ij44 (.clk(clk),.A(search[((8*((17*3)+12+2))-1):(8*((17*3)+12+1))]),.B(current[((8*((16*3)+12+1))-1):(8*((16*3)+12))]),.AD(difference_matrix[3][12]));
me_PE PE_ij45 (.clk(clk),.A(search[((8*((17*3)+13+2))-1):(8*((17*3)+13+1))]),.B(current[((8*((16*3)+13+1))-1):(8*((16*3)+13))]),.AD(difference_matrix[3][13]));
me_PE PE_ij46 (.clk(clk),.A(search[((8*((17*3)+14+2))-1):(8*((17*3)+14+1))]),.B(current[((8*((16*3)+14+1))-1):(8*((16*3)+14))]),.AD(difference_matrix[3][14]));
me_PE PE_ij47 (.clk(clk),.A(search[((8*((17*3)+15+2))-1):(8*((17*3)+15+1))]),.B(current[((8*((16*3)+15+1))-1):(8*((16*3)+15))]),.AD(difference_matrix[3][15]));

me_PE PE_ij64 (.clk(clk),.A(search[((8*((17*4)+0 +2))-1):(8*((17*4)+0 +1))]),.B(current[((8*((16*4)+0 +1))-1):(8*((16*4)+0 ))]),.AD(difference_matrix[4][0 ]));
me_PE PE_ij49 (.clk(clk),.A(search[((8*((17*4)+1 +2))-1):(8*((17*4)+1 +1))]),.B(current[((8*((16*4)+1 +1))-1):(8*((16*4)+1 ))]),.AD(difference_matrix[4][1 ]));
me_PE PE_ij50 (.clk(clk),.A(search[((8*((17*4)+2 +2))-1):(8*((17*4)+2 +1))]),.B(current[((8*((16*4)+2 +1))-1):(8*((16*4)+2 ))]),.AD(difference_matrix[4][2 ]));
me_PE PE_ij51 (.clk(clk),.A(search[((8*((17*4)+3 +2))-1):(8*((17*4)+3 +1))]),.B(current[((8*((16*4)+3 +1))-1):(8*((16*4)+3 ))]),.AD(difference_matrix[4][3 ]));
me_PE PE_ij52 (.clk(clk),.A(search[((8*((17*4)+4 +2))-1):(8*((17*4)+4 +1))]),.B(current[((8*((16*4)+4 +1))-1):(8*((16*4)+4 ))]),.AD(difference_matrix[4][4 ]));
me_PE PE_ij53 (.clk(clk),.A(search[((8*((17*4)+5 +2))-1):(8*((17*4)+5 +1))]),.B(current[((8*((16*4)+5 +1))-1):(8*((16*4)+5 ))]),.AD(difference_matrix[4][5 ]));
me_PE PE_ij54 (.clk(clk),.A(search[((8*((17*4)+6 +2))-1):(8*((17*4)+6 +1))]),.B(current[((8*((16*4)+6 +1))-1):(8*((16*4)+6 ))]),.AD(difference_matrix[4][6 ]));
me_PE PE_ij55 (.clk(clk),.A(search[((8*((17*4)+7 +2))-1):(8*((17*4)+7 +1))]),.B(current[((8*((16*4)+7 +1))-1):(8*((16*4)+7 ))]),.AD(difference_matrix[4][7 ]));
me_PE PE_ij56 (.clk(clk),.A(search[((8*((17*4)+8 +2))-1):(8*((17*4)+8 +1))]),.B(current[((8*((16*4)+8 +1))-1):(8*((16*4)+8 ))]),.AD(difference_matrix[4][8 ]));
me_PE PE_ij57 (.clk(clk),.A(search[((8*((17*4)+9 +2))-1):(8*((17*4)+9 +1))]),.B(current[((8*((16*4)+9 +1))-1):(8*((16*4)+9 ))]),.AD(difference_matrix[4][9 ]));
me_PE PE_ij58 (.clk(clk),.A(search[((8*((17*4)+10+2))-1):(8*((17*4)+10+1))]),.B(current[((8*((16*4)+10+1))-1):(8*((16*4)+10))]),.AD(difference_matrix[4][10]));
me_PE PE_ij59 (.clk(clk),.A(search[((8*((17*4)+11+2))-1):(8*((17*4)+11+1))]),.B(current[((8*((16*4)+11+1))-1):(8*((16*4)+11))]),.AD(difference_matrix[4][11]));
me_PE PE_ij60 (.clk(clk),.A(search[((8*((17*4)+12+2))-1):(8*((17*4)+12+1))]),.B(current[((8*((16*4)+12+1))-1):(8*((16*4)+12))]),.AD(difference_matrix[4][12]));
me_PE PE_ij61 (.clk(clk),.A(search[((8*((17*4)+13+2))-1):(8*((17*4)+13+1))]),.B(current[((8*((16*4)+13+1))-1):(8*((16*4)+13))]),.AD(difference_matrix[4][13]));
me_PE PE_ij62 (.clk(clk),.A(search[((8*((17*4)+14+2))-1):(8*((17*4)+14+1))]),.B(current[((8*((16*4)+14+1))-1):(8*((16*4)+14))]),.AD(difference_matrix[4][14]));
me_PE PE_ij63 (.clk(clk),.A(search[((8*((17*4)+15+2))-1):(8*((17*4)+15+1))]),.B(current[((8*((16*4)+15+1))-1):(8*((16*4)+15))]),.AD(difference_matrix[4][15]));


me_PE PE_ij80 (.clk(clk),.A(search[((8*((17*5)+0 +2))-1):(8*((17*5)+0 +1))]),.B(current[((8*((16*5)+0 +1))-1):(8*((16*5)+0 ))]),.AD(difference_matrix[5][0 ]));
me_PE PE_ij65 (.clk(clk),.A(search[((8*((17*5)+1 +2))-1):(8*((17*5)+1 +1))]),.B(current[((8*((16*5)+1 +1))-1):(8*((16*5)+1 ))]),.AD(difference_matrix[5][1 ]));
me_PE PE_ij66 (.clk(clk),.A(search[((8*((17*5)+2 +2))-1):(8*((17*5)+2 +1))]),.B(current[((8*((16*5)+2 +1))-1):(8*((16*5)+2 ))]),.AD(difference_matrix[5][2 ]));
me_PE PE_ij67 (.clk(clk),.A(search[((8*((17*5)+3 +2))-1):(8*((17*5)+3 +1))]),.B(current[((8*((16*5)+3 +1))-1):(8*((16*5)+3 ))]),.AD(difference_matrix[5][3 ]));
me_PE PE_ij68 (.clk(clk),.A(search[((8*((17*5)+4 +2))-1):(8*((17*5)+4 +1))]),.B(current[((8*((16*5)+4 +1))-1):(8*((16*5)+4 ))]),.AD(difference_matrix[5][4 ]));
me_PE PE_ij69 (.clk(clk),.A(search[((8*((17*5)+5 +2))-1):(8*((17*5)+5 +1))]),.B(current[((8*((16*5)+5 +1))-1):(8*((16*5)+5 ))]),.AD(difference_matrix[5][5 ]));
me_PE PE_ij70 (.clk(clk),.A(search[((8*((17*5)+6 +2))-1):(8*((17*5)+6 +1))]),.B(current[((8*((16*5)+6 +1))-1):(8*((16*5)+6 ))]),.AD(difference_matrix[5][6 ]));
me_PE PE_ij71 (.clk(clk),.A(search[((8*((17*5)+7 +2))-1):(8*((17*5)+7 +1))]),.B(current[((8*((16*5)+7 +1))-1):(8*((16*5)+7 ))]),.AD(difference_matrix[5][7 ]));
me_PE PE_ij72 (.clk(clk),.A(search[((8*((17*5)+8 +2))-1):(8*((17*5)+8 +1))]),.B(current[((8*((16*5)+8 +1))-1):(8*((16*5)+8 ))]),.AD(difference_matrix[5][8 ]));
me_PE PE_ij73 (.clk(clk),.A(search[((8*((17*5)+9 +2))-1):(8*((17*5)+9 +1))]),.B(current[((8*((16*5)+9 +1))-1):(8*((16*5)+9 ))]),.AD(difference_matrix[5][9 ]));
me_PE PE_ij74 (.clk(clk),.A(search[((8*((17*5)+10+2))-1):(8*((17*5)+10+1))]),.B(current[((8*((16*5)+10+1))-1):(8*((16*5)+10))]),.AD(difference_matrix[5][10]));
me_PE PE_ij75 (.clk(clk),.A(search[((8*((17*5)+11+2))-1):(8*((17*5)+11+1))]),.B(current[((8*((16*5)+11+1))-1):(8*((16*5)+11))]),.AD(difference_matrix[5][11]));
me_PE PE_ij76 (.clk(clk),.A(search[((8*((17*5)+12+2))-1):(8*((17*5)+12+1))]),.B(current[((8*((16*5)+12+1))-1):(8*((16*5)+12))]),.AD(difference_matrix[5][12]));
me_PE PE_ij77 (.clk(clk),.A(search[((8*((17*5)+13+2))-1):(8*((17*5)+13+1))]),.B(current[((8*((16*5)+13+1))-1):(8*((16*5)+13))]),.AD(difference_matrix[5][13]));
me_PE PE_ij78 (.clk(clk),.A(search[((8*((17*5)+14+2))-1):(8*((17*5)+14+1))]),.B(current[((8*((16*5)+14+1))-1):(8*((16*5)+14))]),.AD(difference_matrix[5][14]));
me_PE PE_ij79 (.clk(clk),.A(search[((8*((17*5)+15+2))-1):(8*((17*5)+15+1))]),.B(current[((8*((16*5)+15+1))-1):(8*((16*5)+15))]),.AD(difference_matrix[5][15]));


me_PE PE_ij96 (.clk(clk),.A(search[((8*((17*6)+0 +2))-1):(8*((17*6)+0 +1))]),.B(current[((8*((16*6)+0 +1))-1):(8*((16*6)+0 ))]),.AD(difference_matrix[6][0 ]));
me_PE PE_ij81 (.clk(clk),.A(search[((8*((17*6)+1 +2))-1):(8*((17*6)+1 +1))]),.B(current[((8*((16*6)+1 +1))-1):(8*((16*6)+1 ))]),.AD(difference_matrix[6][1 ]));
me_PE PE_ij82 (.clk(clk),.A(search[((8*((17*6)+2 +2))-1):(8*((17*6)+2 +1))]),.B(current[((8*((16*6)+2 +1))-1):(8*((16*6)+2 ))]),.AD(difference_matrix[6][2 ]));
me_PE PE_ij83 (.clk(clk),.A(search[((8*((17*6)+3 +2))-1):(8*((17*6)+3 +1))]),.B(current[((8*((16*6)+3 +1))-1):(8*((16*6)+3 ))]),.AD(difference_matrix[6][3 ]));
me_PE PE_ij84 (.clk(clk),.A(search[((8*((17*6)+4 +2))-1):(8*((17*6)+4 +1))]),.B(current[((8*((16*6)+4 +1))-1):(8*((16*6)+4 ))]),.AD(difference_matrix[6][4 ]));
me_PE PE_ij85 (.clk(clk),.A(search[((8*((17*6)+5 +2))-1):(8*((17*6)+5 +1))]),.B(current[((8*((16*6)+5 +1))-1):(8*((16*6)+5 ))]),.AD(difference_matrix[6][5 ]));
me_PE PE_ij86 (.clk(clk),.A(search[((8*((17*6)+6 +2))-1):(8*((17*6)+6 +1))]),.B(current[((8*((16*6)+6 +1))-1):(8*((16*6)+6 ))]),.AD(difference_matrix[6][6 ]));
me_PE PE_ij87 (.clk(clk),.A(search[((8*((17*6)+7 +2))-1):(8*((17*6)+7 +1))]),.B(current[((8*((16*6)+7 +1))-1):(8*((16*6)+7 ))]),.AD(difference_matrix[6][7 ]));
me_PE PE_ij88 (.clk(clk),.A(search[((8*((17*6)+8 +2))-1):(8*((17*6)+8 +1))]),.B(current[((8*((16*6)+8 +1))-1):(8*((16*6)+8 ))]),.AD(difference_matrix[6][8 ]));
me_PE PE_ij89 (.clk(clk),.A(search[((8*((17*6)+9 +2))-1):(8*((17*6)+9 +1))]),.B(current[((8*((16*6)+9 +1))-1):(8*((16*6)+9 ))]),.AD(difference_matrix[6][9 ]));
me_PE PE_ij90 (.clk(clk),.A(search[((8*((17*6)+10+2))-1):(8*((17*6)+10+1))]),.B(current[((8*((16*6)+10+1))-1):(8*((16*6)+10))]),.AD(difference_matrix[6][10]));
me_PE PE_ij91 (.clk(clk),.A(search[((8*((17*6)+11+2))-1):(8*((17*6)+11+1))]),.B(current[((8*((16*6)+11+1))-1):(8*((16*6)+11))]),.AD(difference_matrix[6][11]));
me_PE PE_ij92 (.clk(clk),.A(search[((8*((17*6)+12+2))-1):(8*((17*6)+12+1))]),.B(current[((8*((16*6)+12+1))-1):(8*((16*6)+12))]),.AD(difference_matrix[6][12]));
me_PE PE_ij93 (.clk(clk),.A(search[((8*((17*6)+13+2))-1):(8*((17*6)+13+1))]),.B(current[((8*((16*6)+13+1))-1):(8*((16*6)+13))]),.AD(difference_matrix[6][13]));
me_PE PE_ij94 (.clk(clk),.A(search[((8*((17*6)+14+2))-1):(8*((17*6)+14+1))]),.B(current[((8*((16*6)+14+1))-1):(8*((16*6)+14))]),.AD(difference_matrix[6][14]));
me_PE PE_ij95 (.clk(clk),.A(search[((8*((17*6)+15+2))-1):(8*((17*6)+15+1))]),.B(current[((8*((16*6)+15+1))-1):(8*((16*6)+15))]),.AD(difference_matrix[6][15]));

me_PE PE_ij112 (.clk(clk),.A(search[((8*((17*7)+0 +2))-1):(8*((17*7)+0 +1))]),.B(current[((8*((16*7)+0 +1))-1):(8*((16*7)+0 ))]),.AD(difference_matrix[7][0 ]));
me_PE PE_ij97 (.clk(clk),.A(search[((8*((17*7)+1 +2))-1):(8*((17*7)+1 +1))]),.B(current[((8*((16*7)+1 +1))-1):(8*((16*7)+1 ))]),.AD(difference_matrix[7][1 ]));
me_PE PE_ij98 (.clk(clk),.A(search[((8*((17*7)+2 +2))-1):(8*((17*7)+2 +1))]),.B(current[((8*((16*7)+2 +1))-1):(8*((16*7)+2 ))]),.AD(difference_matrix[7][2 ]));
me_PE PE_ij99 (.clk(clk),.A(search[((8*((17*7)+3 +2))-1):(8*((17*7)+3 +1))]),.B(current[((8*((16*7)+3 +1))-1):(8*((16*7)+3 ))]),.AD(difference_matrix[7][3 ]));
me_PE PE_ij100 (.clk(clk),.A(search[((8*((17*7)+4 +2))-1):(8*((17*7)+4 +1))]),.B(current[((8*((16*7)+4 +1))-1):(8*((16*7)+4 ))]),.AD(difference_matrix[7][4 ]));
me_PE PE_ij101 (.clk(clk),.A(search[((8*((17*7)+5 +2))-1):(8*((17*7)+5 +1))]),.B(current[((8*((16*7)+5 +1))-1):(8*((16*7)+5 ))]),.AD(difference_matrix[7][5 ]));
me_PE PE_ij102 (.clk(clk),.A(search[((8*((17*7)+6 +2))-1):(8*((17*7)+6 +1))]),.B(current[((8*((16*7)+6 +1))-1):(8*((16*7)+6 ))]),.AD(difference_matrix[7][6 ]));
me_PE PE_ij103 (.clk(clk),.A(search[((8*((17*7)+7 +2))-1):(8*((17*7)+7 +1))]),.B(current[((8*((16*7)+7 +1))-1):(8*((16*7)+7 ))]),.AD(difference_matrix[7][7 ]));
me_PE PE_ij104 (.clk(clk),.A(search[((8*((17*7)+8 +2))-1):(8*((17*7)+8 +1))]),.B(current[((8*((16*7)+8 +1))-1):(8*((16*7)+8 ))]),.AD(difference_matrix[7][8 ]));
me_PE PE_ij105 (.clk(clk),.A(search[((8*((17*7)+9 +2))-1):(8*((17*7)+9 +1))]),.B(current[((8*((16*7)+9 +1))-1):(8*((16*7)+9 ))]),.AD(difference_matrix[7][9 ]));
me_PE PE_ij106 (.clk(clk),.A(search[((8*((17*7)+10+2))-1):(8*((17*7)+10+1))]),.B(current[((8*((16*7)+10+1))-1):(8*((16*7)+10))]),.AD(difference_matrix[7][10]));
me_PE PE_ij107 (.clk(clk),.A(search[((8*((17*7)+11+2))-1):(8*((17*7)+11+1))]),.B(current[((8*((16*7)+11+1))-1):(8*((16*7)+11))]),.AD(difference_matrix[7][11]));
me_PE PE_ij108 (.clk(clk),.A(search[((8*((17*7)+12+2))-1):(8*((17*7)+12+1))]),.B(current[((8*((16*7)+12+1))-1):(8*((16*7)+12))]),.AD(difference_matrix[7][12]));
me_PE PE_ij109 (.clk(clk),.A(search[((8*((17*7)+13+2))-1):(8*((17*7)+13+1))]),.B(current[((8*((16*7)+13+1))-1):(8*((16*7)+13))]),.AD(difference_matrix[7][13]));
me_PE PE_ij110 (.clk(clk),.A(search[((8*((17*7)+14+2))-1):(8*((17*7)+14+1))]),.B(current[((8*((16*7)+14+1))-1):(8*((16*7)+14))]),.AD(difference_matrix[7][14]));
me_PE PE_ij111 (.clk(clk),.A(search[((8*((17*7)+15+2))-1):(8*((17*7)+15+1))]),.B(current[((8*((16*7)+15+1))-1):(8*((16*7)+15))]),.AD(difference_matrix[7][15]));


me_PE PE_ij128 (.clk(clk),.A(search[((8*((17*8)+0 +2))-1):(8*((17*8)+0 +1))]),.B(current[((8*((16*8)+0 +1))-1):(8*((16*8)+0 ))]),.AD(difference_matrix[8][0 ]));
me_PE PE_ij113 (.clk(clk),.A(search[((8*((17*8)+1 +2))-1):(8*((17*8)+1 +1))]),.B(current[((8*((16*8)+1 +1))-1):(8*((16*8)+1 ))]),.AD(difference_matrix[8][1 ]));
me_PE PE_ij114 (.clk(clk),.A(search[((8*((17*8)+2 +2))-1):(8*((17*8)+2 +1))]),.B(current[((8*((16*8)+2 +1))-1):(8*((16*8)+2 ))]),.AD(difference_matrix[8][2 ]));
me_PE PE_ij115 (.clk(clk),.A(search[((8*((17*8)+3 +2))-1):(8*((17*8)+3 +1))]),.B(current[((8*((16*8)+3 +1))-1):(8*((16*8)+3 ))]),.AD(difference_matrix[8][3 ]));
me_PE PE_ij116 (.clk(clk),.A(search[((8*((17*8)+4 +2))-1):(8*((17*8)+4 +1))]),.B(current[((8*((16*8)+4 +1))-1):(8*((16*8)+4 ))]),.AD(difference_matrix[8][4 ]));
me_PE PE_ij117 (.clk(clk),.A(search[((8*((17*8)+5 +2))-1):(8*((17*8)+5 +1))]),.B(current[((8*((16*8)+5 +1))-1):(8*((16*8)+5 ))]),.AD(difference_matrix[8][5 ]));
me_PE PE_ij118 (.clk(clk),.A(search[((8*((17*8)+6 +2))-1):(8*((17*8)+6 +1))]),.B(current[((8*((16*8)+6 +1))-1):(8*((16*8)+6 ))]),.AD(difference_matrix[8][6 ]));
me_PE PE_ij119 (.clk(clk),.A(search[((8*((17*8)+7 +2))-1):(8*((17*8)+7 +1))]),.B(current[((8*((16*8)+7 +1))-1):(8*((16*8)+7 ))]),.AD(difference_matrix[8][7 ]));
me_PE PE_ij120 (.clk(clk),.A(search[((8*((17*8)+8 +2))-1):(8*((17*8)+8 +1))]),.B(current[((8*((16*8)+8 +1))-1):(8*((16*8)+8 ))]),.AD(difference_matrix[8][8 ]));
me_PE PE_ij121 (.clk(clk),.A(search[((8*((17*8)+9 +2))-1):(8*((17*8)+9 +1))]),.B(current[((8*((16*8)+9 +1))-1):(8*((16*8)+9 ))]),.AD(difference_matrix[8][9 ]));
me_PE PE_ij122 (.clk(clk),.A(search[((8*((17*8)+10+2))-1):(8*((17*8)+10+1))]),.B(current[((8*((16*8)+10+1))-1):(8*((16*8)+10))]),.AD(difference_matrix[8][10]));
me_PE PE_ij123 (.clk(clk),.A(search[((8*((17*8)+11+2))-1):(8*((17*8)+11+1))]),.B(current[((8*((16*8)+11+1))-1):(8*((16*8)+11))]),.AD(difference_matrix[8][11]));
me_PE PE_ij124 (.clk(clk),.A(search[((8*((17*8)+12+2))-1):(8*((17*8)+12+1))]),.B(current[((8*((16*8)+12+1))-1):(8*((16*8)+12))]),.AD(difference_matrix[8][12]));
me_PE PE_ij125 (.clk(clk),.A(search[((8*((17*8)+13+2))-1):(8*((17*8)+13+1))]),.B(current[((8*((16*8)+13+1))-1):(8*((16*8)+13))]),.AD(difference_matrix[8][13]));
me_PE PE_ij126 (.clk(clk),.A(search[((8*((17*8)+14+2))-1):(8*((17*8)+14+1))]),.B(current[((8*((16*8)+14+1))-1):(8*((16*8)+14))]),.AD(difference_matrix[8][14]));
me_PE PE_ij127 (.clk(clk),.A(search[((8*((17*8)+15+2))-1):(8*((17*8)+15+1))]),.B(current[((8*((16*8)+15+1))-1):(8*((16*8)+15))]),.AD(difference_matrix[8][15]));

me_PE PE_ij144 (.clk(clk),.A(search[((8*((17*9)+0 +2))-1):(8*((17*9)+0 +1))]),.B(current[((8*((16*9)+0 +1))-1):(8*((16*9)+0 ))]),.AD(difference_matrix[9][0 ]));
me_PE PE_ij129 (.clk(clk),.A(search[((8*((17*9)+1 +2))-1):(8*((17*9)+1 +1))]),.B(current[((8*((16*9)+1 +1))-1):(8*((16*9)+1 ))]),.AD(difference_matrix[9][1 ]));
me_PE PE_ij130 (.clk(clk),.A(search[((8*((17*9)+2 +2))-1):(8*((17*9)+2 +1))]),.B(current[((8*((16*9)+2 +1))-1):(8*((16*9)+2 ))]),.AD(difference_matrix[9][2 ]));
me_PE PE_ij131 (.clk(clk),.A(search[((8*((17*9)+3 +2))-1):(8*((17*9)+3 +1))]),.B(current[((8*((16*9)+3 +1))-1):(8*((16*9)+3 ))]),.AD(difference_matrix[9][3 ]));
me_PE PE_ij132 (.clk(clk),.A(search[((8*((17*9)+4 +2))-1):(8*((17*9)+4 +1))]),.B(current[((8*((16*9)+4 +1))-1):(8*((16*9)+4 ))]),.AD(difference_matrix[9][4 ]));
me_PE PE_ij133 (.clk(clk),.A(search[((8*((17*9)+5 +2))-1):(8*((17*9)+5 +1))]),.B(current[((8*((16*9)+5 +1))-1):(8*((16*9)+5 ))]),.AD(difference_matrix[9][5 ]));
me_PE PE_ij134 (.clk(clk),.A(search[((8*((17*9)+6 +2))-1):(8*((17*9)+6 +1))]),.B(current[((8*((16*9)+6 +1))-1):(8*((16*9)+6 ))]),.AD(difference_matrix[9][6 ]));
me_PE PE_ij135 (.clk(clk),.A(search[((8*((17*9)+7 +2))-1):(8*((17*9)+7 +1))]),.B(current[((8*((16*9)+7 +1))-1):(8*((16*9)+7 ))]),.AD(difference_matrix[9][7 ]));
me_PE PE_ij136 (.clk(clk),.A(search[((8*((17*9)+8 +2))-1):(8*((17*9)+8 +1))]),.B(current[((8*((16*9)+8 +1))-1):(8*((16*9)+8 ))]),.AD(difference_matrix[9][8 ]));
me_PE PE_ij137 (.clk(clk),.A(search[((8*((17*9)+9 +2))-1):(8*((17*9)+9 +1))]),.B(current[((8*((16*9)+9 +1))-1):(8*((16*9)+9 ))]),.AD(difference_matrix[9][9 ]));
me_PE PE_ij138 (.clk(clk),.A(search[((8*((17*9)+10+2))-1):(8*((17*9)+10+1))]),.B(current[((8*((16*9)+10+1))-1):(8*((16*9)+10))]),.AD(difference_matrix[9][10]));
me_PE PE_ij139 (.clk(clk),.A(search[((8*((17*9)+11+2))-1):(8*((17*9)+11+1))]),.B(current[((8*((16*9)+11+1))-1):(8*((16*9)+11))]),.AD(difference_matrix[9][11]));
me_PE PE_ij140 (.clk(clk),.A(search[((8*((17*9)+12+2))-1):(8*((17*9)+12+1))]),.B(current[((8*((16*9)+12+1))-1):(8*((16*9)+12))]),.AD(difference_matrix[9][12]));
me_PE PE_ij141 (.clk(clk),.A(search[((8*((17*9)+13+2))-1):(8*((17*9)+13+1))]),.B(current[((8*((16*9)+13+1))-1):(8*((16*9)+13))]),.AD(difference_matrix[9][13]));
me_PE PE_ij142 (.clk(clk),.A(search[((8*((17*9)+14+2))-1):(8*((17*9)+14+1))]),.B(current[((8*((16*9)+14+1))-1):(8*((16*9)+14))]),.AD(difference_matrix[9][14]));
me_PE PE_ij143 (.clk(clk),.A(search[((8*((17*9)+15+2))-1):(8*((17*9)+15+1))]),.B(current[((8*((16*9)+15+1))-1):(8*((16*9)+15))]),.AD(difference_matrix[9][15]));

me_PE PE_ij160 (.clk(clk),.A(search[((8*((17*10)+0 +2))-1):(8*((17*10)+0 +1))]),.B(current[((8*((16*10)+0 +1))-1):(8*((16*10)+0 ))]),.AD(difference_matrix[10][0 ]));
me_PE PE_ij145 (.clk(clk),.A(search[((8*((17*10)+1 +2))-1):(8*((17*10)+1 +1))]),.B(current[((8*((16*10)+1 +1))-1):(8*((16*10)+1 ))]),.AD(difference_matrix[10][1 ]));
me_PE PE_ij146 (.clk(clk),.A(search[((8*((17*10)+2 +2))-1):(8*((17*10)+2 +1))]),.B(current[((8*((16*10)+2 +1))-1):(8*((16*10)+2 ))]),.AD(difference_matrix[10][2 ]));
me_PE PE_ij147 (.clk(clk),.A(search[((8*((17*10)+3 +2))-1):(8*((17*10)+3 +1))]),.B(current[((8*((16*10)+3 +1))-1):(8*((16*10)+3 ))]),.AD(difference_matrix[10][3 ]));
me_PE PE_ij148 (.clk(clk),.A(search[((8*((17*10)+4 +2))-1):(8*((17*10)+4 +1))]),.B(current[((8*((16*10)+4 +1))-1):(8*((16*10)+4 ))]),.AD(difference_matrix[10][4 ]));
me_PE PE_ij149 (.clk(clk),.A(search[((8*((17*10)+5 +2))-1):(8*((17*10)+5 +1))]),.B(current[((8*((16*10)+5 +1))-1):(8*((16*10)+5 ))]),.AD(difference_matrix[10][5 ]));
me_PE PE_ij150 (.clk(clk),.A(search[((8*((17*10)+6 +2))-1):(8*((17*10)+6 +1))]),.B(current[((8*((16*10)+6 +1))-1):(8*((16*10)+6 ))]),.AD(difference_matrix[10][6 ]));
me_PE PE_ij151 (.clk(clk),.A(search[((8*((17*10)+7 +2))-1):(8*((17*10)+7 +1))]),.B(current[((8*((16*10)+7 +1))-1):(8*((16*10)+7 ))]),.AD(difference_matrix[10][7 ]));
me_PE PE_ij152 (.clk(clk),.A(search[((8*((17*10)+8 +2))-1):(8*((17*10)+8 +1))]),.B(current[((8*((16*10)+8 +1))-1):(8*((16*10)+8 ))]),.AD(difference_matrix[10][8 ]));
me_PE PE_ij153 (.clk(clk),.A(search[((8*((17*10)+9 +2))-1):(8*((17*10)+9 +1))]),.B(current[((8*((16*10)+9 +1))-1):(8*((16*10)+9 ))]),.AD(difference_matrix[10][9 ]));
me_PE PE_ij154 (.clk(clk),.A(search[((8*((17*10)+10+2))-1):(8*((17*10)+10+1))]),.B(current[((8*((16*10)+10+1))-1):(8*((16*10)+10))]),.AD(difference_matrix[10][10]));
me_PE PE_ij155 (.clk(clk),.A(search[((8*((17*10)+11+2))-1):(8*((17*10)+11+1))]),.B(current[((8*((16*10)+11+1))-1):(8*((16*10)+11))]),.AD(difference_matrix[10][11]));
me_PE PE_ij156 (.clk(clk),.A(search[((8*((17*10)+12+2))-1):(8*((17*10)+12+1))]),.B(current[((8*((16*10)+12+1))-1):(8*((16*10)+12))]),.AD(difference_matrix[10][12]));
me_PE PE_ij157 (.clk(clk),.A(search[((8*((17*10)+13+2))-1):(8*((17*10)+13+1))]),.B(current[((8*((16*10)+13+1))-1):(8*((16*10)+13))]),.AD(difference_matrix[10][13]));
me_PE PE_ij158 (.clk(clk),.A(search[((8*((17*10)+14+2))-1):(8*((17*10)+14+1))]),.B(current[((8*((16*10)+14+1))-1):(8*((16*10)+14))]),.AD(difference_matrix[10][14]));
me_PE PE_ij159 (.clk(clk),.A(search[((8*((17*10)+15+2))-1):(8*((17*10)+15+1))]),.B(current[((8*((16*10)+15+1))-1):(8*((16*10)+15))]),.AD(difference_matrix[10][15]));
           
me_PE PE_ij176 (.clk(clk),.A(search[((8*((17*11)+0 +2))-1):(8*((17*11)+0 +1))]),.B(current[((8*((16*11)+0 +1))-1):(8*((16*11)+0 ))]),.AD(difference_matrix[11][0 ]));
me_PE PE_ij161 (.clk(clk),.A(search[((8*((17*11)+1 +2))-1):(8*((17*11)+1 +1))]),.B(current[((8*((16*11)+1 +1))-1):(8*((16*11)+1 ))]),.AD(difference_matrix[11][1 ]));
me_PE PE_ij162 (.clk(clk),.A(search[((8*((17*11)+2 +2))-1):(8*((17*11)+2 +1))]),.B(current[((8*((16*11)+2 +1))-1):(8*((16*11)+2 ))]),.AD(difference_matrix[11][2 ]));
me_PE PE_ij163 (.clk(clk),.A(search[((8*((17*11)+3 +2))-1):(8*((17*11)+3 +1))]),.B(current[((8*((16*11)+3 +1))-1):(8*((16*11)+3 ))]),.AD(difference_matrix[11][3 ]));
me_PE PE_ij164 (.clk(clk),.A(search[((8*((17*11)+4 +2))-1):(8*((17*11)+4 +1))]),.B(current[((8*((16*11)+4 +1))-1):(8*((16*11)+4 ))]),.AD(difference_matrix[11][4 ]));
me_PE PE_ij165 (.clk(clk),.A(search[((8*((17*11)+5 +2))-1):(8*((17*11)+5 +1))]),.B(current[((8*((16*11)+5 +1))-1):(8*((16*11)+5 ))]),.AD(difference_matrix[11][5 ]));
me_PE PE_ij166 (.clk(clk),.A(search[((8*((17*11)+6 +2))-1):(8*((17*11)+6 +1))]),.B(current[((8*((16*11)+6 +1))-1):(8*((16*11)+6 ))]),.AD(difference_matrix[11][6 ]));
me_PE PE_ij167 (.clk(clk),.A(search[((8*((17*11)+7 +2))-1):(8*((17*11)+7 +1))]),.B(current[((8*((16*11)+7 +1))-1):(8*((16*11)+7 ))]),.AD(difference_matrix[11][7 ]));
me_PE PE_ij168 (.clk(clk),.A(search[((8*((17*11)+8 +2))-1):(8*((17*11)+8 +1))]),.B(current[((8*((16*11)+8 +1))-1):(8*((16*11)+8 ))]),.AD(difference_matrix[11][8 ]));
me_PE PE_ij169 (.clk(clk),.A(search[((8*((17*11)+9 +2))-1):(8*((17*11)+9 +1))]),.B(current[((8*((16*11)+9 +1))-1):(8*((16*11)+9 ))]),.AD(difference_matrix[11][9 ]));
me_PE PE_ij170 (.clk(clk),.A(search[((8*((17*11)+10+2))-1):(8*((17*11)+10+1))]),.B(current[((8*((16*11)+10+1))-1):(8*((16*11)+10))]),.AD(difference_matrix[11][10]));
me_PE PE_ij171 (.clk(clk),.A(search[((8*((17*11)+11+2))-1):(8*((17*11)+11+1))]),.B(current[((8*((16*11)+11+1))-1):(8*((16*11)+11))]),.AD(difference_matrix[11][11]));
me_PE PE_ij172 (.clk(clk),.A(search[((8*((17*11)+12+2))-1):(8*((17*11)+12+1))]),.B(current[((8*((16*11)+12+1))-1):(8*((16*11)+12))]),.AD(difference_matrix[11][12]));
me_PE PE_ij173 (.clk(clk),.A(search[((8*((17*11)+13+2))-1):(8*((17*11)+13+1))]),.B(current[((8*((16*11)+13+1))-1):(8*((16*11)+13))]),.AD(difference_matrix[11][13]));
me_PE PE_ij174 (.clk(clk),.A(search[((8*((17*11)+14+2))-1):(8*((17*11)+14+1))]),.B(current[((8*((16*11)+14+1))-1):(8*((16*11)+14))]),.AD(difference_matrix[11][14]));
me_PE PE_ij175 (.clk(clk),.A(search[((8*((17*11)+15+2))-1):(8*((17*11)+15+1))]),.B(current[((8*((16*11)+15+1))-1):(8*((16*11)+15))]),.AD(difference_matrix[11][15]));

me_PE PE_ij192 (.clk(clk),.A(search[((8*((17*12)+0 +2))-1):(8*((17*12)+0 +1))]),.B(current[((8*((16*12)+0 +1))-1):(8*((16*12)+0 ))]),.AD(difference_matrix[12][0 ]));
me_PE PE_ij177 (.clk(clk),.A(search[((8*((17*12)+1 +2))-1):(8*((17*12)+1 +1))]),.B(current[((8*((16*12)+1 +1))-1):(8*((16*12)+1 ))]),.AD(difference_matrix[12][1 ]));
me_PE PE_ij178 (.clk(clk),.A(search[((8*((17*12)+2 +2))-1):(8*((17*12)+2 +1))]),.B(current[((8*((16*12)+2 +1))-1):(8*((16*12)+2 ))]),.AD(difference_matrix[12][2 ]));
me_PE PE_ij179 (.clk(clk),.A(search[((8*((17*12)+3 +2))-1):(8*((17*12)+3 +1))]),.B(current[((8*((16*12)+3 +1))-1):(8*((16*12)+3 ))]),.AD(difference_matrix[12][3 ]));
me_PE PE_ij180 (.clk(clk),.A(search[((8*((17*12)+4 +2))-1):(8*((17*12)+4 +1))]),.B(current[((8*((16*12)+4 +1))-1):(8*((16*12)+4 ))]),.AD(difference_matrix[12][4 ]));
me_PE PE_ij181 (.clk(clk),.A(search[((8*((17*12)+5 +2))-1):(8*((17*12)+5 +1))]),.B(current[((8*((16*12)+5 +1))-1):(8*((16*12)+5 ))]),.AD(difference_matrix[12][5 ]));
me_PE PE_ij182 (.clk(clk),.A(search[((8*((17*12)+6 +2))-1):(8*((17*12)+6 +1))]),.B(current[((8*((16*12)+6 +1))-1):(8*((16*12)+6 ))]),.AD(difference_matrix[12][6 ]));
me_PE PE_ij183 (.clk(clk),.A(search[((8*((17*12)+7 +2))-1):(8*((17*12)+7 +1))]),.B(current[((8*((16*12)+7 +1))-1):(8*((16*12)+7 ))]),.AD(difference_matrix[12][7 ]));
me_PE PE_ij184 (.clk(clk),.A(search[((8*((17*12)+8 +2))-1):(8*((17*12)+8 +1))]),.B(current[((8*((16*12)+8 +1))-1):(8*((16*12)+8 ))]),.AD(difference_matrix[12][8 ]));
me_PE PE_ij185 (.clk(clk),.A(search[((8*((17*12)+9 +2))-1):(8*((17*12)+9 +1))]),.B(current[((8*((16*12)+9 +1))-1):(8*((16*12)+9 ))]),.AD(difference_matrix[12][9 ]));
me_PE PE_ij186 (.clk(clk),.A(search[((8*((17*12)+10+2))-1):(8*((17*12)+10+1))]),.B(current[((8*((16*12)+10+1))-1):(8*((16*12)+10))]),.AD(difference_matrix[12][10]));
me_PE PE_ij187 (.clk(clk),.A(search[((8*((17*12)+11+2))-1):(8*((17*12)+11+1))]),.B(current[((8*((16*12)+11+1))-1):(8*((16*12)+11))]),.AD(difference_matrix[12][11]));
me_PE PE_ij188 (.clk(clk),.A(search[((8*((17*12)+12+2))-1):(8*((17*12)+12+1))]),.B(current[((8*((16*12)+12+1))-1):(8*((16*12)+12))]),.AD(difference_matrix[12][12]));
me_PE PE_ij189 (.clk(clk),.A(search[((8*((17*12)+13+2))-1):(8*((17*12)+13+1))]),.B(current[((8*((16*12)+13+1))-1):(8*((16*12)+13))]),.AD(difference_matrix[12][13]));
me_PE PE_ij190 (.clk(clk),.A(search[((8*((17*12)+14+2))-1):(8*((17*12)+14+1))]),.B(current[((8*((16*12)+14+1))-1):(8*((16*12)+14))]),.AD(difference_matrix[12][14]));
me_PE PE_ij191 (.clk(clk),.A(search[((8*((17*12)+15+2))-1):(8*((17*12)+15+1))]),.B(current[((8*((16*12)+15+1))-1):(8*((16*12)+15))]),.AD(difference_matrix[12][15]));

me_PE PE_ij208 (.clk(clk),.A(search[((8*((17*13)+0 +2))-1):(8*((17*13)+0 +1))]),.B(current[((8*((16*13)+0 +1))-1):(8*((16*13)+0 ))]),.AD(difference_matrix[13][0 ]));
me_PE PE_ij193 (.clk(clk),.A(search[((8*((17*13)+1 +2))-1):(8*((17*13)+1 +1))]),.B(current[((8*((16*13)+1 +1))-1):(8*((16*13)+1 ))]),.AD(difference_matrix[13][1 ]));
me_PE PE_ij194 (.clk(clk),.A(search[((8*((17*13)+2 +2))-1):(8*((17*13)+2 +1))]),.B(current[((8*((16*13)+2 +1))-1):(8*((16*13)+2 ))]),.AD(difference_matrix[13][2 ]));
me_PE PE_ij195 (.clk(clk),.A(search[((8*((17*13)+3 +2))-1):(8*((17*13)+3 +1))]),.B(current[((8*((16*13)+3 +1))-1):(8*((16*13)+3 ))]),.AD(difference_matrix[13][3 ]));
me_PE PE_ij196 (.clk(clk),.A(search[((8*((17*13)+4 +2))-1):(8*((17*13)+4 +1))]),.B(current[((8*((16*13)+4 +1))-1):(8*((16*13)+4 ))]),.AD(difference_matrix[13][4 ]));
me_PE PE_ij197 (.clk(clk),.A(search[((8*((17*13)+5 +2))-1):(8*((17*13)+5 +1))]),.B(current[((8*((16*13)+5 +1))-1):(8*((16*13)+5 ))]),.AD(difference_matrix[13][5 ]));
me_PE PE_ij198 (.clk(clk),.A(search[((8*((17*13)+6 +2))-1):(8*((17*13)+6 +1))]),.B(current[((8*((16*13)+6 +1))-1):(8*((16*13)+6 ))]),.AD(difference_matrix[13][6 ]));
me_PE PE_ij199 (.clk(clk),.A(search[((8*((17*13)+7 +2))-1):(8*((17*13)+7 +1))]),.B(current[((8*((16*13)+7 +1))-1):(8*((16*13)+7 ))]),.AD(difference_matrix[13][7 ]));
me_PE PE_ij200 (.clk(clk),.A(search[((8*((17*13)+8 +2))-1):(8*((17*13)+8 +1))]),.B(current[((8*((16*13)+8 +1))-1):(8*((16*13)+8 ))]),.AD(difference_matrix[13][8 ]));
me_PE PE_ij201 (.clk(clk),.A(search[((8*((17*13)+9 +2))-1):(8*((17*13)+9 +1))]),.B(current[((8*((16*13)+9 +1))-1):(8*((16*13)+9 ))]),.AD(difference_matrix[13][9 ]));
me_PE PE_ij202 (.clk(clk),.A(search[((8*((17*13)+10+2))-1):(8*((17*13)+10+1))]),.B(current[((8*((16*13)+10+1))-1):(8*((16*13)+10))]),.AD(difference_matrix[13][10]));
me_PE PE_ij203 (.clk(clk),.A(search[((8*((17*13)+11+2))-1):(8*((17*13)+11+1))]),.B(current[((8*((16*13)+11+1))-1):(8*((16*13)+11))]),.AD(difference_matrix[13][11]));
me_PE PE_ij204 (.clk(clk),.A(search[((8*((17*13)+12+2))-1):(8*((17*13)+12+1))]),.B(current[((8*((16*13)+12+1))-1):(8*((16*13)+12))]),.AD(difference_matrix[13][12]));
me_PE PE_ij205 (.clk(clk),.A(search[((8*((17*13)+13+2))-1):(8*((17*13)+13+1))]),.B(current[((8*((16*13)+13+1))-1):(8*((16*13)+13))]),.AD(difference_matrix[13][13]));
me_PE PE_ij206 (.clk(clk),.A(search[((8*((17*13)+14+2))-1):(8*((17*13)+14+1))]),.B(current[((8*((16*13)+14+1))-1):(8*((16*13)+14))]),.AD(difference_matrix[13][14]));
me_PE PE_ij207 (.clk(clk),.A(search[((8*((17*13)+15+2))-1):(8*((17*13)+15+1))]),.B(current[((8*((16*13)+15+1))-1):(8*((16*13)+15))]),.AD(difference_matrix[13][15]));

me_PE PE_ij224 (.clk(clk),.A(search[((8*((17*14)+0 +2))-1):(8*((17*14)+0 +1))]),.B(current[((8*((16*14)+0 +1))-1):(8*((16*14)+0 ))]),.AD(difference_matrix[14][0 ]));
me_PE PE_ij209 (.clk(clk),.A(search[((8*((17*14)+1 +2))-1):(8*((17*14)+1 +1))]),.B(current[((8*((16*14)+1 +1))-1):(8*((16*14)+1 ))]),.AD(difference_matrix[14][1 ]));
me_PE PE_ij210 (.clk(clk),.A(search[((8*((17*14)+2 +2))-1):(8*((17*14)+2 +1))]),.B(current[((8*((16*14)+2 +1))-1):(8*((16*14)+2 ))]),.AD(difference_matrix[14][2 ]));
me_PE PE_ij211 (.clk(clk),.A(search[((8*((17*14)+3 +2))-1):(8*((17*14)+3 +1))]),.B(current[((8*((16*14)+3 +1))-1):(8*((16*14)+3 ))]),.AD(difference_matrix[14][3 ]));
me_PE PE_ij212 (.clk(clk),.A(search[((8*((17*14)+4 +2))-1):(8*((17*14)+4 +1))]),.B(current[((8*((16*14)+4 +1))-1):(8*((16*14)+4 ))]),.AD(difference_matrix[14][4 ]));
me_PE PE_ij213 (.clk(clk),.A(search[((8*((17*14)+5 +2))-1):(8*((17*14)+5 +1))]),.B(current[((8*((16*14)+5 +1))-1):(8*((16*14)+5 ))]),.AD(difference_matrix[14][5 ]));
me_PE PE_ij214 (.clk(clk),.A(search[((8*((17*14)+6 +2))-1):(8*((17*14)+6 +1))]),.B(current[((8*((16*14)+6 +1))-1):(8*((16*14)+6 ))]),.AD(difference_matrix[14][6 ]));
me_PE PE_ij215 (.clk(clk),.A(search[((8*((17*14)+7 +2))-1):(8*((17*14)+7 +1))]),.B(current[((8*((16*14)+7 +1))-1):(8*((16*14)+7 ))]),.AD(difference_matrix[14][7 ]));
me_PE PE_ij216 (.clk(clk),.A(search[((8*((17*14)+8 +2))-1):(8*((17*14)+8 +1))]),.B(current[((8*((16*14)+8 +1))-1):(8*((16*14)+8 ))]),.AD(difference_matrix[14][8 ]));
me_PE PE_ij217 (.clk(clk),.A(search[((8*((17*14)+9 +2))-1):(8*((17*14)+9 +1))]),.B(current[((8*((16*14)+9 +1))-1):(8*((16*14)+9 ))]),.AD(difference_matrix[14][9 ]));
me_PE PE_ij218 (.clk(clk),.A(search[((8*((17*14)+10+2))-1):(8*((17*14)+10+1))]),.B(current[((8*((16*14)+10+1))-1):(8*((16*14)+10))]),.AD(difference_matrix[14][10]));
me_PE PE_ij219 (.clk(clk),.A(search[((8*((17*14)+11+2))-1):(8*((17*14)+11+1))]),.B(current[((8*((16*14)+11+1))-1):(8*((16*14)+11))]),.AD(difference_matrix[14][11]));
me_PE PE_ij220 (.clk(clk),.A(search[((8*((17*14)+12+2))-1):(8*((17*14)+12+1))]),.B(current[((8*((16*14)+12+1))-1):(8*((16*14)+12))]),.AD(difference_matrix[14][12]));
me_PE PE_ij221 (.clk(clk),.A(search[((8*((17*14)+13+2))-1):(8*((17*14)+13+1))]),.B(current[((8*((16*14)+13+1))-1):(8*((16*14)+13))]),.AD(difference_matrix[14][13]));
me_PE PE_ij222 (.clk(clk),.A(search[((8*((17*14)+14+2))-1):(8*((17*14)+14+1))]),.B(current[((8*((16*14)+14+1))-1):(8*((16*14)+14))]),.AD(difference_matrix[14][14]));
me_PE PE_ij223 (.clk(clk),.A(search[((8*((17*14)+15+2))-1):(8*((17*14)+15+1))]),.B(current[((8*((16*14)+15+1))-1):(8*((16*14)+15))]),.AD(difference_matrix[14][15]));

me_PE PE_ij240 (.clk(clk),.A(search[((8*((17*15)+0 +2))-1):(8*((17*15)+0 +1))]),.B(current[((8*((16*15)+0 +1))-1):(8*((16*15)+0 ))]),.AD(difference_matrix[15][0 ]));
me_PE PE_ij225 (.clk(clk),.A(search[((8*((17*15)+1 +2))-1):(8*((17*15)+1 +1))]),.B(current[((8*((16*15)+1 +1))-1):(8*((16*15)+1 ))]),.AD(difference_matrix[15][1 ]));
me_PE PE_ij226 (.clk(clk),.A(search[((8*((17*15)+2 +2))-1):(8*((17*15)+2 +1))]),.B(current[((8*((16*15)+2 +1))-1):(8*((16*15)+2 ))]),.AD(difference_matrix[15][2 ]));
me_PE PE_ij227 (.clk(clk),.A(search[((8*((17*15)+3 +2))-1):(8*((17*15)+3 +1))]),.B(current[((8*((16*15)+3 +1))-1):(8*((16*15)+3 ))]),.AD(difference_matrix[15][3 ]));
me_PE PE_ij228 (.clk(clk),.A(search[((8*((17*15)+4 +2))-1):(8*((17*15)+4 +1))]),.B(current[((8*((16*15)+4 +1))-1):(8*((16*15)+4 ))]),.AD(difference_matrix[15][4 ]));
me_PE PE_ij229 (.clk(clk),.A(search[((8*((17*15)+5 +2))-1):(8*((17*15)+5 +1))]),.B(current[((8*((16*15)+5 +1))-1):(8*((16*15)+5 ))]),.AD(difference_matrix[15][5 ]));
me_PE PE_ij230 (.clk(clk),.A(search[((8*((17*15)+6 +2))-1):(8*((17*15)+6 +1))]),.B(current[((8*((16*15)+6 +1))-1):(8*((16*15)+6 ))]),.AD(difference_matrix[15][6 ]));
me_PE PE_ij231 (.clk(clk),.A(search[((8*((17*15)+7 +2))-1):(8*((17*15)+7 +1))]),.B(current[((8*((16*15)+7 +1))-1):(8*((16*15)+7 ))]),.AD(difference_matrix[15][7 ]));
me_PE PE_ij232 (.clk(clk),.A(search[((8*((17*15)+8 +2))-1):(8*((17*15)+8 +1))]),.B(current[((8*((16*15)+8 +1))-1):(8*((16*15)+8 ))]),.AD(difference_matrix[15][8 ]));
me_PE PE_ij233 (.clk(clk),.A(search[((8*((17*15)+9 +2))-1):(8*((17*15)+9 +1))]),.B(current[((8*((16*15)+9 +1))-1):(8*((16*15)+9 ))]),.AD(difference_matrix[15][9 ]));
me_PE PE_ij234 (.clk(clk),.A(search[((8*((17*15)+10+2))-1):(8*((17*15)+10+1))]),.B(current[((8*((16*15)+10+1))-1):(8*((16*15)+10))]),.AD(difference_matrix[15][10]));
me_PE PE_ij235 (.clk(clk),.A(search[((8*((17*15)+11+2))-1):(8*((17*15)+11+1))]),.B(current[((8*((16*15)+11+1))-1):(8*((16*15)+11))]),.AD(difference_matrix[15][11]));
me_PE PE_ij236 (.clk(clk),.A(search[((8*((17*15)+12+2))-1):(8*((17*15)+12+1))]),.B(current[((8*((16*15)+12+1))-1):(8*((16*15)+12))]),.AD(difference_matrix[15][12]));
me_PE PE_ij237 (.clk(clk),.A(search[((8*((17*15)+13+2))-1):(8*((17*15)+13+1))]),.B(current[((8*((16*15)+13+1))-1):(8*((16*15)+13))]),.AD(difference_matrix[15][13]));
me_PE PE_ij238 (.clk(clk),.A(search[((8*((17*15)+14+2))-1):(8*((17*15)+14+1))]),.B(current[((8*((16*15)+14+1))-1):(8*((16*15)+14))]),.AD(difference_matrix[15][14]));
me_PE PE_ij239 (.clk(clk),.A(search[((8*((17*15)+15+2))-1):(8*((17*15)+15+1))]),.B(current[((8*((16*15)+15+1))-1):(8*((16*15)+15))]),.AD(difference_matrix[15][15]));

	
	always @ (posedge clk)
	begin 
		add01	<=	(difference_matrix [0][0][7:0] + difference_matrix [0][1][7:0]) + (difference_matrix [0][2][7:0] + difference_matrix [0][3][7:0]);
		add02	<=	(difference_matrix [0][4][7:0] + difference_matrix [0][5][7:0]) + (difference_matrix [0][6][7:0] + difference_matrix [0][7][7:0]);
		add03	<=	(difference_matrix [0][8][7:0] + difference_matrix [0][9][7:0]) + (difference_matrix [0][10][7:0] + difference_matrix [0][11][7:0]);
		add04	<=	(difference_matrix [0][12][7:0] + difference_matrix [0][13][7:0]) + (difference_matrix [0][14][7:0] + difference_matrix [0][15][7:0]);
		add05	<=	(difference_matrix [1][0][7:0] + difference_matrix [1][1][7:0]) + (difference_matrix [1][2][7:0] + difference_matrix [1][3][7:0]);
		add06	<=	(difference_matrix [1][4][7:0] + difference_matrix [1][5][7:0]) + (difference_matrix [1][6][7:0] + difference_matrix [1][7][7:0]);
		add07	<=	(difference_matrix [1][8][7:0] + difference_matrix [1][9][7:0]) + (difference_matrix [1][10][7:0] + difference_matrix [1][11][7:0]);
		add08	<=	(difference_matrix [1][12][7:0] + difference_matrix [1][13][7:0]) + (difference_matrix [1][14][7:0] + difference_matrix [1][15][7:0]);
		add09	<=	(difference_matrix [2][0][7:0] + difference_matrix [2][1][7:0]) + (difference_matrix [2][2][7:0] + difference_matrix [2][3][7:0]);
		add10	<=	(difference_matrix [2][4][7:0] + difference_matrix [2][5][7:0]) + (difference_matrix [2][6][7:0] + difference_matrix [2][7][7:0]);
		add11	<=	(difference_matrix [2][8][7:0] + difference_matrix [2][9][7:0]) + (difference_matrix [2][10][7:0] + difference_matrix [2][11][7:0]);
		add12	<=	(difference_matrix [2][12][7:0] + difference_matrix [2][13][7:0]) + (difference_matrix [2][14][7:0] + difference_matrix [2][15][7:0]);
		add13	<=	(difference_matrix [3][0][7:0] + difference_matrix [3][1][7:0]) + (difference_matrix [3][2][7:0] + difference_matrix [3][3][7:0]);
		add14	<=	(difference_matrix [3][4][7:0] + difference_matrix [3][5][7:0]) + (difference_matrix [3][6][7:0] + difference_matrix [3][7][7:0]);
		add15	<=	(difference_matrix [3][8][7:0] + difference_matrix [3][9][7:0]) + (difference_matrix [3][10][7:0] + difference_matrix [3][11][7:0]);
		add16	<=	(difference_matrix [3][12][7:0] + difference_matrix [3][13][7:0]) + (difference_matrix [3][14][7:0] + difference_matrix [3][15][7:0]);
		add17	<=	(difference_matrix [4][0][7:0] + difference_matrix [4][1][7:0]) + (difference_matrix [4][2][7:0] + difference_matrix [4][3][7:0]);
		add18	<=	(difference_matrix [4][4][7:0] + difference_matrix [4][5][7:0]) + (difference_matrix [4][6][7:0] + difference_matrix [4][7][7:0]);
		add19	<=	(difference_matrix [4][8][7:0] + difference_matrix [4][9][7:0]) + (difference_matrix [4][10][7:0] + difference_matrix [4][11][7:0]);
		add20	<=	(difference_matrix [4][12][7:0] + difference_matrix [4][13][7:0]) + (difference_matrix [4][14][7:0] + difference_matrix [4][15][7:0]);
		add21	<=	(difference_matrix [5][0][7:0] + difference_matrix [5][1][7:0]) + (difference_matrix [5][2][7:0] + difference_matrix [5][3][7:0]);
		add22	<=	(difference_matrix [5][4][7:0] + difference_matrix [5][5][7:0]) + (difference_matrix [5][6][7:0] + difference_matrix [5][7][7:0]);
		add23	<=	(difference_matrix [5][8][7:0] + difference_matrix [5][9][7:0]) + (difference_matrix [5][10][7:0] + difference_matrix [5][11][7:0]);
		add24	<=	(difference_matrix [5][12][7:0] + difference_matrix [5][13][7:0]) + (difference_matrix [5][14][7:0] + difference_matrix [5][15][7:0]);
		add25	<=	(difference_matrix [6][0][7:0] + difference_matrix [6][1][7:0]) + (difference_matrix [6][2][7:0] + difference_matrix [6][3][7:0]);
		add26	<=	(difference_matrix [6][4][7:0] + difference_matrix [6][5][7:0]) + (difference_matrix [6][6][7:0] + difference_matrix [6][7][7:0]);
		add27	<=	(difference_matrix [6][8][7:0] + difference_matrix [6][9][7:0]) + (difference_matrix [6][10][7:0] + difference_matrix [6][11][7:0]);
		add28	<=	(difference_matrix [6][12][7:0] + difference_matrix [6][13][7:0]) + (difference_matrix [6][14][7:0] + difference_matrix [6][15][7:0]);
		add29	<=	(difference_matrix [7][0][7:0] + difference_matrix [7][1][7:0]) + (difference_matrix [7][2][7:0] + difference_matrix [7][3][7:0]);
		add30	<=	(difference_matrix [7][4][7:0] + difference_matrix [7][5][7:0]) + (difference_matrix [7][6][7:0] + difference_matrix [7][7][7:0]);
		add31	<=	(difference_matrix [7][8][7:0] + difference_matrix [7][9][7:0]) + (difference_matrix [7][10][7:0] + difference_matrix [7][11][7:0]);
		add32	<=	(difference_matrix [7][12][7:0] + difference_matrix [7][13][7:0]) + (difference_matrix [7][14][7:0] + difference_matrix [7][15][7:0]);
		add33	<=	(difference_matrix [8][0][7:0] + difference_matrix [8][1][7:0]) + (difference_matrix [8][2][7:0] + difference_matrix [8][3][7:0]);
		add34	<=	(difference_matrix [8][4][7:0] + difference_matrix [8][5][7:0]) + (difference_matrix [8][6][7:0] + difference_matrix [8][7][7:0]);
		add35	<=	(difference_matrix [8][8][7:0] + difference_matrix [8][9][7:0]) + (difference_matrix [8][10][7:0] + difference_matrix [8][11][7:0]);
		add36	<=	(difference_matrix [8][12][7:0] + difference_matrix [8][13][7:0]) + (difference_matrix [8][14][7:0] + difference_matrix [8][15][7:0]);
		add37	<=	(difference_matrix [9][0][7:0] + difference_matrix [9][1][7:0]) + (difference_matrix [9][2][7:0] + difference_matrix [9][3][7:0]);
		add38	<=	(difference_matrix [9][4][7:0] + difference_matrix [9][5][7:0]) + (difference_matrix [9][6][7:0] + difference_matrix [9][7][7:0]);
		add39	<=	(difference_matrix [9][8][7:0] + difference_matrix [9][9][7:0]) + (difference_matrix [9][10][7:0] + difference_matrix [9][11][7:0]);
		add40	<=	(difference_matrix [9][12][7:0] + difference_matrix [9][13][7:0]) + (difference_matrix [9][14][7:0] + difference_matrix [9][15][7:0]);
		add41	<=	(difference_matrix [10][0][7:0] + difference_matrix [10][1][7:0]) + (difference_matrix [10][2][7:0] + difference_matrix [10][3][7:0]);
		add42	<=	(difference_matrix [10][4][7:0] + difference_matrix [10][5][7:0]) + (difference_matrix [10][6][7:0] + difference_matrix [10][7][7:0]);
		add43	<=	(difference_matrix [10][8][7:0] + difference_matrix [10][9][7:0]) + (difference_matrix [10][10][7:0] + difference_matrix [10][11][7:0]);
		add44	<=	(difference_matrix [10][12][7:0] + difference_matrix [10][13][7:0]) + (difference_matrix [10][14][7:0] + difference_matrix [10][15][7:0]);
		add45	<=	(difference_matrix [11][0][7:0] + difference_matrix [11][1][7:0]) + (difference_matrix [11][2][7:0] + difference_matrix [11][3][7:0]);
		add46	<=	(difference_matrix [11][4][7:0] + difference_matrix [11][5][7:0]) + (difference_matrix [11][6][7:0] + difference_matrix [11][7][7:0]);
		add47	<=	(difference_matrix [11][8][7:0] + difference_matrix [11][9][7:0]) + (difference_matrix [11][10][7:0] + difference_matrix [11][11][7:0]);
		add48	<=	(difference_matrix [11][12][7:0] + difference_matrix [11][13][7:0]) + (difference_matrix [11][14][7:0] + difference_matrix [11][15][7:0]);
		add49	<=	(difference_matrix [12][0][7:0] + difference_matrix [12][1][7:0]) + (difference_matrix [12][2][7:0] + difference_matrix [12][3][7:0]);
		add50	<=	(difference_matrix [12][4][7:0] + difference_matrix [12][5][7:0]) + (difference_matrix [12][6][7:0] + difference_matrix [12][7][7:0]);
		add51	<=	(difference_matrix [12][8][7:0] + difference_matrix [12][9][7:0]) + (difference_matrix [12][10][7:0] + difference_matrix [12][11][7:0]);
		add52	<=	(difference_matrix [12][12][7:0] + difference_matrix [12][13][7:0]) + (difference_matrix [12][14][7:0] + difference_matrix [12][15][7:0]);
		add53	<=	(difference_matrix [13][0][7:0] + difference_matrix [13][1][7:0]) + (difference_matrix [13][2][7:0] + difference_matrix [13][3][7:0]);
		add54	<=	(difference_matrix [13][4][7:0] + difference_matrix [13][5][7:0]) + (difference_matrix [13][6][7:0] + difference_matrix [13][7][7:0]);
		add55	<=	(difference_matrix [13][8][7:0] + difference_matrix [13][9][7:0]) + (difference_matrix [13][10][7:0] + difference_matrix [13][11][7:0]);
		add56	<=	(difference_matrix [13][12][7:0] + difference_matrix [13][13][7:0]) + (difference_matrix [13][14][7:0] + difference_matrix [13][15][7:0]);
		add57	<=	(difference_matrix [14][0][7:0] + difference_matrix [14][1][7:0]) + (difference_matrix [14][2][7:0] + difference_matrix [14][3][7:0]);
		add58	<=	(difference_matrix [14][4][7:0] + difference_matrix [14][5][7:0]) + (difference_matrix [14][6][7:0] + difference_matrix [14][7][7:0]);
		add59	<=	(difference_matrix [14][8][7:0] + difference_matrix [14][9][7:0]) + (difference_matrix [14][10][7:0] + difference_matrix [14][11][7:0]);
		add60	<=	(difference_matrix [14][12][7:0] + difference_matrix [14][13][7:0]) + (difference_matrix [14][14][7:0] + difference_matrix [14][15][7:0]);
		add61	<=	(difference_matrix [15][0][7:0] + difference_matrix [15][1][7:0]) + (difference_matrix [15][2][7:0] + difference_matrix [15][3][7:0]);
		add62	<=	(difference_matrix [15][4][7:0] + difference_matrix [15][5][7:0]) + (difference_matrix [15][6][7:0] + difference_matrix [15][7][7:0]);
		add63	<=	(difference_matrix [15][8][7:0] + difference_matrix [15][9][7:0]) + (difference_matrix [15][10][7:0] + difference_matrix [15][11][7:0]);
		add64	<=	(difference_matrix [15][12][7:0] + difference_matrix [15][13][7:0]) + (difference_matrix [15][14][7:0] + difference_matrix [15][15][7:0]);
	end
	
	always @ (posedge clk)
	begin
		SAD01 <= (add52 + add56) + (add60 + add64);
		SAD02 <= (add51 + add55) + (add59 + add63);
		SAD03 <= (add50 + add54) + (add58 + add62);
		SAD04 <= (add49 + add53) + (add57 + add61);
		SAD05 <= (add36 + add40) + (add44 + add48);
		SAD06 <= (add35 + add39) + (add43 + add47);
		SAD07 <= (add34 + add38) + (add42 + add46);
		SAD08 <= (add33 + add37) + (add41 + add45);
		SAD09 <= (add20 + add24) + (add28 + add32);
		SAD10 <= (add19 + add23) + (add27 + add31);
		SAD11 <= (add18 + add22) + (add26 + add30);
		SAD12 <= (add17 + add21) + (add25 + add29);
		SAD13 <= (add04 + add08) + (add12 + add16);
		SAD14 <= (add03 + add07) + (add11 + add15);
		SAD15 <= (add02 + add06) + (add10 + add14);
		SAD16 <= (add01 + add05) + (add09 + add13);
	end
endmodule
